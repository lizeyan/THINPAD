----------------------------------------------------------------------------------
-- Company: Concept Computer Corporation
-- Engineer: LXH, LZY, YST
-- 
-- Create Date:    11:15:22 11/18/2016 
-- Design Name: 
-- Module Name:    ControlUnit - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;

entity ControlUnit is
    Port ( 
           -- IF generate
           ExDigitsOp : out STD_LOGIC_VECTOR(2 downto 0); --���䵽ExtendModule
           ExSignOp : out STD_LOGIC;
           -- ID
           AluOp : out STD_LOGIC_VECTOR(3 downto 0); -- ���浽ID_RF
           AMuxOp : out STD_LOGIC_VECTOR(3 downto 0); --
           BMuxOp : out STD_LOGIC_VECTOR(2 downto 0); --
           DirOp : out STD_LOGIC_VECTOR(2 downto 0); -- ���䵽DirectionModule
           IDPCOp : out STD_LOGIC_VECTOR(1 downto 0); 
           
           RegWrbOp : out STD_LOGIC_VECTOR(1 downto 0); -- �Ĵ���д�����ݵ�ѡ�� -- ���浽ID_RF
           RXTOp : out STD_LOGIC_VECTOR(2 downto 0);
           SWSrc : out STD_LOGIC; -- 0 rx, 1 ry --���浽ID_RF
           RamRWOp : out STD_LOGIC; -- 0 read, 1 write --���浽ID_RF
           BTBOP : out STD_LOGIC; -- is jumping ins(1) or not(0)
                -- ENABLE  complex
           EXE_RFOp : out STD_LOGIC_VECTOR(1 downto 0);
           ID_RFOp : out STD_LOGIC_VECTOR(1 downto 0);
           IF_RFOp : out STD_LOGIC_VECTOR(1 downto 0);
           MEM_RFOp : out STD_LOGIC_VECTOR(1 downto 0);
           PC_RFOp : out STD_LOGIC_VECTOR(2 downto 0);
           
			  -- ��IF�θոմ��ڴ���ȡ�������ʵ�ָ��
           PC_RF_PC: in STD_LOGIC_VECTOR (15 downto 0);
           IF_Ins : in STD_LOGIC_VECTOR(15 downto 0);
           
           IF_RF_OP : in STD_LOGIC_VECTOR(4 downto 0);
           IF_RF_ST: in STD_LOGIC_VECTOR (15 downto 0); -- IF�μĴ����б���ģ�ָ������ݡ���Ϊ�е�ָ����Ҫ�ж�funct�ֶ�
           IDPC: in STD_LOGIC_VECTOR (15 downto 0); -- IDPCRXT������IDPC
           ID_RF_OP : in STD_LOGIC_VECTOR(4 downto 0); 
           ID_RF_Rd : in STD_LOGIC_VECTOR(3 downto 0);
           EXE_RF_OP : in STD_LOGIC_VECTOR(4 downto 0);
           EXE_RF_Rd : in STD_LOGIC_VECTOR(3 downto 0);
           EXE_Fout : in STD_LOGIC_VECTOR (15 downto 0); -- ALU�ļ�ʱ���
           MEM_RF_OP : in STD_LOGIC_VECTOR(4 downto 0);
           MEM_RF_Rd : in STD_LOGIC_VECTOR(3 downto 0)
           );
end ControlUnit;

architecture Behavioral of ControlUnit is
	---------------------------------------------------------------------------------------------
    function last_lw_rd (signal x: STD_LOGIC_VECTOR (3 downto 0)) 
		return boolean is
	 begin
		return ((ID_RF_RD = x) and (ID_RF_OP = "10010" or ID_RF_OP = "10011"));
	 end last_lw_rd;
	 -----------------------------------------------------------------------------------------------
	 -- 111�Ƿ�����ʾNone
	 signal PC_SRC_IF, PC_SRC_ID, PC_SRC_EXE, PC_SRC_MEM, PC_SRC_WB: STD_LOGIC_VECTOR (2 downto 0) := "000";
begin
	-- ����MEM_RFOP
	mem_rfop <= "00";
	
	-- ����EXE_RFOP
	exe_rfop <= "00";

    -- generate btbop signal
    process(if_rf_st)
        variable op = if_rf_st(15 downto 11);
    begin
        if(op="00010" or op="00100" or op="00101") -- b, beqz, bnez
            btbop <= '1';
        elsif(if_rf_st(15 downto 8)="01100000")  -- bteqz
            btbop <= '1';
        elsif(op="11101" and if_rf_st="00000") -- jr
            btbop <= '1';
        else
            btbop <= '0';
        end if;
    end process;
    
	--���������ж�������࣬������д��һ��process���棬̫������дһ�����
	-- ������ܲ��㣬���Բ𿪳�����process�ֱ����
	-- ����ID_RFOP
	-- ����IF_RFOP
	process (if_rf_st, pc_rf_pc, idpc, id_rf_op, id_rf_rd, exe_rf_op, exe_rf_rd)
		variable target_failed : boolean := false; --��תָ���Ԥ��ʧ��
		variable last_lw_rd, last_last_lw_rd, last_rd : boolean := false; --�������ݳ�ͻ
		variable written_st: boolean := false; --����֮����swָ����д���ָ��ĵ�ַ
		--------------------------------------------------------------------------------------------------
		procedure data_conflict (x: in std_logic_vector(3 downto 0);
--														signal id_rf_rd, exe_rf_rd: in std_logic_vector (3 downto 0);
--														signal id_rf_op, exe_rf_op: in std_logic_vector (4 downto 0);
													  last_rd, last_lw_rd, last_last_lw_rd: out boolean) is
		begin
			last_rd := id_rf_rd = x;
			last_lw_rd := (id_rf_rd = x) and (id_rf_op = "10011" or id_rf_op = "10010");
			last_last_lw_rd := (exe_rf_op = "10011" or exe_rf_op = "10010") and exe_rf_rd = x;
		end data_conflict;
		procedure data_conflict (x, y: in std_logic_vector(3 downto 0);
--														signal id_rf_rd, exe_rf_rd: in std_logic_vector (3 downto 0);
--														signal id_rf_op, exe_rf_op: in std_logic_vector (4 downto 0);
													  last_rd, last_lw_rd, last_last_lw_rd: out boolean) is
		begin
			last_rd := id_rf_rd = x or id_rf_rd = y;
			last_lw_rd := (id_rf_rd = x or id_rf_rd = y) and (id_rf_op = "10011" or id_rf_op = "10010");
			last_last_lw_rd := (exe_rf_op = "10011" or exe_rf_op = "10010") and (exe_rf_rd = x or exe_rf_rd = y);
		end data_conflict;
		procedure normal_ins(last_rd, last_lw_rd, last_last_lw_rd, written_st, target_failed: in boolean) is
		begin
				if written_st then
					if_rfop <= "11";
					id_rfop <= "11";
				elsif last_lw_rd then
					if_rfop <= "10";
					id_rfop <= "11";
				else
					if_rfop <= "00";
					id_rfop <= "00";
				end if;
		end normal_ins;
		procedure branch_ins(last_rd, last_lw_rd, last_last_lw_rd, written_st, target_failed: in boolean) is
		begin
			if written_st or (target_failed and not (last_rd or last_last_lw_rd)) then
				if_rfop <= "11";
				id_rfop <= "11";
			elsif last_rd or last_last_lw_rd then
				if_rfop <= "10";
				id_rfop <= "11";
			else
				if_rfop <= "00";
				id_rfop <= "00";
			end if;
		end branch_ins;
	begin
		target_failed := idpc /= pc_rf_pc;
		---------------------------------------------------------------------------------
		written_st := (id_rf_op = "11011" or id_rf_op = "11010") and exe_fout = pc_rf_pc;
		---------------------------------------------------------------------------------
		case if_rf_st(15 downto 11) is
			when "01001" => -- addiu
				data_conflict (x => '0' & if_rf_st(10 downto 8), last_rd => last_rd, last_lw_rd => last_lw_rd, last_last_lw_rd => last_last_lw_rd);
				normal_ins (last_rd => last_rd, last_lw_rd => last_lw_rd, last_last_lw_rd => last_last_lw_rd, written_st => written_st, target_failed => target_failed);
			when "01000" => -- addiu3
				data_conflict (x => '0' & if_rf_st(10 downto 8), last_rd => last_rd, last_lw_rd => last_lw_rd, last_last_lw_rd => last_last_lw_rd);
				normal_ins (last_rd => last_rd, last_lw_rd => last_lw_rd, last_last_lw_rd => last_last_lw_rd, written_st => written_st, target_failed => target_failed);
			when "01100" => 
				case if_rf_st (10 downto 8) is
					when "011" => -- addsp
						data_conflict (x => "1001", last_rd => last_rd, last_lw_rd => last_lw_rd, last_last_lw_rd => last_last_lw_rd);
						normal_ins (last_rd => last_rd, last_lw_rd => last_lw_rd, last_last_lw_rd => last_last_lw_rd, written_st => written_st, target_failed => target_failed);
					when "000" => --btnez
						data_conflict (x => "1010", last_rd => last_rd, last_lw_rd => last_lw_rd, last_last_lw_rd => last_last_lw_rd);
						branch_ins (last_rd => last_rd, last_lw_rd => last_lw_rd, last_last_lw_rd => last_last_lw_rd, written_st => written_st, target_failed => target_failed);
					when "100" => --mtsp
							data_conflict (x => '0' & if_rf_st(7 downto 5), last_rd => last_rd, last_lw_rd => last_lw_rd, last_last_lw_rd => last_last_lw_rd);
						normal_ins (last_rd => last_rd, last_lw_rd => last_lw_rd, last_last_lw_rd => last_last_lw_rd, written_st => written_st, target_failed => target_failed);
					when others =>
						if_rfop <= "00";
				end case;
			when "00000" => --addsp3
				data_conflict (x => "1001", last_rd => last_rd, last_lw_rd => last_lw_rd, last_last_lw_rd => last_last_lw_rd);
				normal_ins (last_rd => last_rd, last_lw_rd => last_lw_rd, last_last_lw_rd => last_last_lw_rd, written_st => written_st, target_failed => target_failed);
			when "00010" => -- b
				normal_ins (last_rd => last_rd, last_lw_rd => last_lw_rd, last_last_lw_rd => last_last_lw_rd, written_st => written_st, target_failed => target_failed);
			when "00100" => -- beqz
				data_conflict (x => '0' & if_rf_st(10 downto 8), last_rd => last_rd, last_lw_rd => last_lw_rd, last_last_lw_rd => last_last_lw_rd);
				branch_ins (last_rd => last_rd, last_lw_rd => last_lw_rd, last_last_lw_rd => last_last_lw_rd, written_st => written_st, target_failed => target_failed);
			when "00101" => -- bnez
				data_conflict (x => '0' & if_rf_st(10 downto 8), last_rd => last_rd, last_lw_rd => last_lw_rd, last_last_lw_rd => last_last_lw_rd);
				branch_ins (last_rd => last_rd, last_lw_rd => last_lw_rd, last_last_lw_rd => last_last_lw_rd, written_st => written_st, target_failed => target_failed);
			when "01110" => -- cmpi
				data_conflict (x => '0' & if_rf_st(10 downto 8), last_rd => last_rd, last_lw_rd => last_lw_rd, last_last_lw_rd => last_last_lw_rd);
				normal_ins (last_rd => last_rd, last_lw_rd => last_lw_rd, last_last_lw_rd => last_last_lw_rd, written_st => written_st, target_failed => target_failed);
			when "01101" => -- li
				normal_ins (last_rd => last_rd, last_lw_rd => last_lw_rd, last_last_lw_rd => last_last_lw_rd, written_st => written_st, target_failed => target_failed);
			when "10011" => -- lw
				data_conflict (x => '0' & if_rf_st(10 downto 8), last_rd => last_rd, last_lw_rd => last_lw_rd, last_last_lw_rd => last_last_lw_rd);
				normal_ins (last_rd => last_rd, last_lw_rd => last_lw_rd, last_last_lw_rd => last_last_lw_rd, written_st => written_st, target_failed => target_failed);
			when "10010" => -- lw_sp
				data_conflict (x => "1001", last_rd => last_rd, last_lw_rd => last_lw_rd, last_last_lw_rd => last_last_lw_rd);
				normal_ins (last_rd => last_rd, last_lw_rd => last_lw_rd, last_last_lw_rd => last_last_lw_rd, written_st => written_st, target_failed => target_failed);
			when "00110" => -- sll, sra
				case if_rf_st(1 downto 0) is
					when "00" =>
						data_conflict (x => '0' & if_rf_st(7 downto 5), last_rd => last_rd, last_lw_rd => last_lw_rd, last_last_lw_rd => last_last_lw_rd);
					when "11" =>
						data_conflict (x => '0' & if_rf_st(7 downto 5), last_rd => last_rd, last_lw_rd => last_lw_rd, last_last_lw_rd => last_last_lw_rd);
					when others =>
				end case;
				normal_ins (last_rd => last_rd, last_lw_rd => last_lw_rd, last_last_lw_rd => last_last_lw_rd, written_st => written_st, target_failed => target_failed);
			when "01010" => -- slti
				data_conflict (x => '0' & if_rf_st(10 downto 8), y => '0' & if_rf_st(7 downto 5), last_rd => last_rd, last_lw_rd => last_lw_rd, last_last_lw_rd => last_last_lw_rd);
				normal_ins (last_rd => last_rd, last_lw_rd => last_lw_rd, last_last_lw_rd => last_last_lw_rd, written_st => written_st, target_failed => target_failed);
			when "01111" => --move
				data_conflict (x => '0' & if_rf_st(7 downto 5), last_rd => last_rd, last_lw_rd => last_lw_rd, last_last_lw_rd => last_last_lw_rd);
				normal_ins (last_rd => last_rd, last_lw_rd => last_lw_rd, last_last_lw_rd => last_last_lw_rd, written_st => written_st, target_failed => target_failed);
			when "11011" => -- sw
				data_conflict (x => '0' & if_rf_st(10 downto 8), y => '0' & if_rf_st(7 downto 5), last_rd => last_rd, last_lw_rd => last_lw_rd, last_last_lw_rd => last_last_lw_rd);
				normal_ins (last_rd => last_rd, last_lw_rd => last_lw_rd, last_last_lw_rd => last_last_lw_rd, written_st => written_st, target_failed => target_failed);
			when "11010" => -- swsp
				data_conflict (x => '0' & if_rf_st(10 downto 8), y => "1001", last_rd => last_rd, last_lw_rd => last_lw_rd, last_last_lw_rd => last_last_lw_rd);
				normal_ins (last_rd => last_rd, last_lw_rd => last_lw_rd, last_last_lw_rd => last_last_lw_rd, written_st => written_st, target_failed => target_failed);
			when "11100" => 
				case if_rf_st(1 downto 0) is
					when "01" => --addu
						data_conflict (x => '0' & if_rf_st(10 downto 8), y => '0' & if_rf_st(7 downto 5), last_rd => last_rd, last_lw_rd => last_lw_rd, last_last_lw_rd => last_last_lw_rd);
					when "11" => --subu
						data_conflict (x => '0' & if_rf_st(10 downto 8), y => '0' & if_rf_st(7 downto 5), last_rd => last_rd, last_lw_rd => last_lw_rd, last_last_lw_rd => last_last_lw_rd);
					when others =>
				end case;
				normal_ins (last_rd => last_rd, last_lw_rd => last_lw_rd, last_last_lw_rd => last_last_lw_rd, written_st => written_st, target_failed => target_failed);
			when "11101" =>
				case if_rf_st(4 downto 0) is
					when "01100" => -- add
						normal_ins (last_rd => last_rd, last_lw_rd => last_lw_rd, last_last_lw_rd => last_last_lw_rd, written_st => written_st, target_failed => target_failed);
					when "01010" => --cmp
						data_conflict (x => '0' & if_rf_st(10 downto 8), y => '0' & if_rf_st(7 downto 5), last_rd => last_rd, last_lw_rd => last_lw_rd, last_last_lw_rd => last_last_lw_rd);
						normal_ins (last_rd => last_rd, last_lw_rd => last_lw_rd, last_last_lw_rd => last_last_lw_rd, written_st => written_st, target_failed => target_failed);
					when "11101" => --or
						data_conflict (x => '0' & if_rf_st(10 downto 8), y => '0' & if_rf_st(7 downto 5), last_rd => last_rd, last_lw_rd => last_lw_rd, last_last_lw_rd => last_last_lw_rd);
						normal_ins (last_rd => last_rd, last_lw_rd => last_lw_rd, last_last_lw_rd => last_last_lw_rd, written_st => written_st, target_failed => target_failed);
					when "00100" => -- sllv
						data_conflict (x => '0' & if_rf_st(10 downto 8), y => '0' & if_rf_st(7 downto 5), last_rd => last_rd, last_lw_rd => last_lw_rd, last_last_lw_rd => last_last_lw_rd);
						normal_ins (last_rd => last_rd, last_lw_rd => last_lw_rd, last_last_lw_rd => last_last_lw_rd, written_st => written_st, target_failed => target_failed);
					when "00000" => 
						if if_rf_st(7 downto 5) = "0000" then --jr
							data_conflict (x => '0' & if_rf_st(10 downto 8), last_rd => last_rd, last_lw_rd => last_lw_rd, last_last_lw_rd => last_last_lw_rd);
								branch_ins (last_rd => last_rd, last_lw_rd => last_lw_rd, last_last_lw_rd => last_last_lw_rd, written_st => written_st, target_failed => target_failed);
						elsif if_rf_st(7 downto 5) = "0100" then --mfpc
								normal_ins (last_rd => last_rd, last_lw_rd => last_lw_rd, last_last_lw_rd => last_last_lw_rd, written_st => written_st, target_failed => target_failed);
						else
						end if;
					when others =>
				end case;
			when "11110" => --mfih and mtih
				case if_rf_st(0) is
					when '0' => -- mfih
					when '1' => -- mtih
						data_conflict (x => '0' & if_rf_st(10 downto 8), last_rd => last_rd, last_lw_rd => last_lw_rd, last_last_lw_rd => last_last_lw_rd);
					when others =>
				end case;
				normal_ins (last_rd => last_rd, last_lw_rd => last_lw_rd, last_last_lw_rd => last_last_lw_rd, written_st => written_st, target_failed => target_failed);
			when "11111" => --int
				if_rfop <= "00";
				id_rfop <= "00";
			when others =>
				normal_ins (last_rd => last_rd, last_lw_rd => last_lw_rd, last_last_lw_rd => last_last_lw_rd, written_st => written_st, target_failed => target_failed);
		end case;
	end process;

	-- ����RXTOP��Ȼ�󴫸�IDPCRXTʹ�ã�������
	-- ʹ��IF�μĴ����е�ָ���ֶ�
	process (if_rf_st)
		-- 00 x
		-- 10 exe_rf_res
		-- 11 mem_rf_lw
		-- 01 mem_rf_res
		variable x : STD_LOGIC_VECTOR (3 downto 0) := "1111"; --����ָ����Ҫ�ļĴ����ĵ�ַ
	begin
		-- ȷ��������תָ����Ҫ�ļĴ�����ַ
		if if_rf_st(15 downto 11) = "00010" then --b
			x := "1111";
		elsif if_rf_st(15 downto 11) = "00100" then --beqz
			x := '0' & if_rf_st (10 downto 8);
		elsif if_rf_st(15 downto 11) = "00101" then --bnez
			x := '0' & if_rf_st (10 downto 8);
		elsif if_rf_st(15 downto 8) = "01100000" then --bteqz
			x := "1010";
		elsif if_rf_st(15 downto 11) = "11101" and if_rf_st(7 downto 0) = "00000000" then --jr
			x := '0' & if_rf_st (10 downto 8);
		else
			x := "1111";
		end if;
		-- ����б�Ҫȡ�Ĵ�����ֵ
		if x /= "1111" then --�Ͳ鿴֮ǰָ��������ʹ��������·
			if id_rf_rd = x then --�����һ��ָ���ַ��ͬ����Ҫ�ȴ�һ�غϣ���������ѡ���ﲢ���ؼ�
				rxtop <= "000"; -- useless
			else
				if exe_rf_rd = x then --���������ָ���lwָ���ô����ȷ������ǵĻ���������Ҫ�ȴ�һ�غϣ����Բ����ؼ�
					rxtop <= "010";
				else
					if mem_rf_rd = x then
						if mem_rf_op = "10011" or mem_rf_op = "10010" then
							rxtop <= "011";
						else
							rxtop <= "100";
						end if;
					else
						if x = "1010" then
							rxtop <= "001";
						else
							rxtop <= "000";
						end if;
					end if;
				end if;
			end if;
		else --���û��Ҫ
			rxtop <= "111"; --�͸����Ƿ������ź�
		end if;
	end process;
    
	-- ����IDPCOP��Ȼ�󴫸�IDPCRXTʹ�ã�������
	-- ʹ��IF�μĴ����е�ָ���ֶ�
	process (if_rf_st)
	begin
		if if_rf_st(15 downto 11) = "00010" then --b
			idpcop <= "10";
		elsif if_rf_st(15 downto 11) = "00100" then --beqz
			idpcop <= "00";
		elsif if_rf_st(15 downto 11) = "00101" then --bnez
			idpcop <= "01";
		elsif if_rf_st(15 downto 8) = "01100000" then --bteqz
			idpcop <= "00";
		elsif if_rf_st(15 downto 11) = "11101" and if_rf_st(7 downto 0) = "00000000" then --jr
			idpcop <= "11";
		else
			idpcop <= "ZZ";
		end if;
	end process;
	--------------------------------------------------------------------------------------------
	--------------------------------------------------------------------------------------------
	--------------------------------------------------------------------------------------------
	-- ����PC_RFOP
	-- pc_src_if
	-- ����INTӦ�õ��쳣�����ַ����Ķ�Ӧ�õ�Ԥ���ַ
	process (if_ins)
	begin
		if if_ins(15 downto 11) = "11111" then --intָ��
			pc_src_if <= "010";
		else
			pc_src_if <= "000";
		end if;
	end process;
    
    
	-- pc_src_id
	-- ����תָ���PDT
	-- ��תָ��Ƚ�Ŀ���PC_RF_PC����ͬ����PDT���������IDPC
	process (if_rf_st)
	begin
		if idpc = pc_rf_pc then
			pc_src_id <= "000";
		else
			pc_src_id <= "001";
		end if;
	end process;
	-- pc_src_exe
	pc_src_exe <= "111";
	-- pc_src_mem
	pc_src_mem <= "111";
	-- pc_src_wb
	pc_src_wb <= "111";
	--�ۺ�
    -- 000 PDTPC
    -- 001 IDPC
    -- 010 �쳣�����ַ
    -- 011 IF_RF_PC_ORIGIN
    -- 100 ����д
	process (pc_src_if, pc_src_id, pc_src_exe, pc_src_mem, pc_src_wb)
	begin
		if pc_src_wb = "111" then
			if pc_src_mem = "111" then
				if pc_src_exe = "111" then
					if pc_src_id = "111" then
						pc_rfop <= pc_src_if;
					else
						pc_rfop <= pc_src_id;
					end if;
				else
					pc_rfop <= pc_src_exe;
				end if;
			else
				pc_rfop <= pc_src_mem;
			end if;
		else
			pc_rfop <= pc_src_wb;
		end if;
	end process;
	--------------------------------------------------------------------------------------------
	--------------------------------------------------------------------------------------------
	--------------------------------------------------------------------------------------------

	-- ����regwrbop, ��֮����Ҫ���䱣�浽ID_RF
	-- ����ramrwop��֮����Ҫ���䱣�浽ID_RF
	-- ����mem_sw_srcop��֮����Ҫ���䱣�浽ID_RF
	-- ����Ŀ��Ĵ���ѡ��Ŀ����룬֮����Ҫ���䴫�䵽DirectionModule
    --- 000 rx
    --- 001 ry
    --- 011 rz
    --- 010 SP
    --- 110 IH
    --- 100 T
    --- others 1111 ILLEGAL
	-- ����ALU�����룬֮����Ҫ���䱣�浽ID_RF
	-- ʹ��ID�εõ���IF_RD_OP
	process (IF_RF_ST)
		variable op: STD_LOGIC_VECTOR (4 downto 0);
		variable dir: STD_LOGIC_VECTOR (2 downto 0); -- 
	begin
		op := if_rf_st (15 downto 11);
		case op is
            when "01001" => -- addiu
					aluop <= "0000";
					dir := "000";
					regwrbop <= "00";
					ramrwop <= '0';
					swsrc <= '0';
            when "01000" => -- addiu3
					aluop <= "0000";
					dir := "001";
					regwrbop <= "00";
					ramrwop <= '0';
					swsrc <= '0';
            when "01100" => --addsp, bteqz, mtsp
					ramrwop <= '0';
					swsrc <= '0';
					case if_rf_st (10 downto 8) is
						when "011" => -- addsp
							aluop <= "0000";
							dir := "010";
							regwrbop <= "00";
						when "000" => --btnez
							aluop <= "0110";
							dir := "111";
							regwrbop <= "11";
						when "100" => --mtsp
							aluop <= "0011";
							dir := "010";
							regwrbop <= "00";
						when others =>
							aluop <= "1111";
							dir := "111";
							regwrbop <= "11";
					end case;
            when "00000" => --addsp3
					ramrwop <= '0';
					swsrc <= '0';
					aluop <= "0000";
					dir := "000";
					regwrbop <= "00";
            when "00010" => -- b
					ramrwop <= '0';
					swsrc <= '0';
					aluop <= "0000";
					dir := "111";
					regwrbop <= "11";
            when "00100" => -- beqz
					ramrwop <= '0';
					swsrc <= '0';
					aluop <= "0110";
					dir := "111";
					regwrbop <= "11";
            when "00101" => -- bnez
					ramrwop <= '0';
					swsrc <= '0';
					aluop <= "0110";
					dir := "111";
					regwrbop <= "11";
            when "01110" => -- cmpi
					ramrwop <= '0';
					swsrc <= '0';
					aluop <= "0110";
					dir := "100";
					regwrbop <= "10";
            when "01101" => -- li
					ramrwop <= '0';
					swsrc <= '0';
					aluop <= "0011";
					dir := "000";
					regwrbop <= "00";
            when "10011" => -- lw
					ramrwop <= '0';
					swsrc <= '0';
					aluop <= "0000";
					dir := "001";
					regwrbop <= "01";
            when "10010" => -- lw_sp
					ramrwop <= '0';
					swsrc <= '0';
					aluop <= "0000";
					dir := "000";
					regwrbop <= "01";
            when "00110" => 
					ramrwop <= '0';
					swsrc <= '0';
					case if_rf_st(1 downto 0) is
					when "00" => --sll
						aluop <= "0111";
						dir := "000";
						regwrbop <= "00";
					when "11" =>
						aluop <= "0100"; --sra
						dir := "000";
						regwrbop <= "00";
					when others =>
						aluop <= "1111";
						dir := "111";
					end case;
            when "01010" => -- slti
					ramrwop <= '0';
					swsrc <= '0';
					aluop <= "0001";
					dir := "100";
					regwrbop <= "00";
				when "01111" => --move
					ramrwop <= '0';
					swsrc <= '0';
					aluop <= "0011";
					dir := "000";
					regwrbop <= "00";
            when "11011" => -- sw
					aluop <= "0000";
					dir := "111";
					ramrwop <= '1';
					swsrc <= '1';
					regwrbop <= "11";
            when "11010" => -- swsp
					aluop <= "0000";
					dir := "111";
					ramrwop <= '1';
					swsrc <= '0';
					regwrbop <= "11";
				when "11100" => 
					ramrwop <= '0';
					swsrc <= '0';
					case if_rf_st(1 downto 0) is
						when "01" => --addu
							aluop <= "0000";
							dir := "011";
							regwrbop <= "00";
						when "11" => --subu
							aluop <= "0001";
							regwrbop <= "00";
							dir := "011";
						when others =>
							aluop <= "1111";
							dir := "111";
					end case;
				when "11101" =>
					ramrwop <= '0';
					swsrc <= '0';
					case if_rf_st(4 downto 0) is
						when "01100" => -- and
							aluop <= "0011";
							dir := "000";
							regwrbop <= "00";
						when "01010" => --cmp
							aluop <= "0110";
							dir := "100";
							regwrbop <= "10";
						when "11101" => --or
							aluop <= "0010";
							dir := "000";
							regwrbop <= "00";
						when "00100" => -- sllv
							aluop <= "0101";
							dir := "001";
							regwrbop <= "00";
						when "00000" => --mfpc
							aluop <= "0010";
							dir := "000";
							regwrbop <= "00";
						when others =>
							aluop <= "1111";
							dir := "111";
							regwrbop <= "11";
					end case;
				when "11110" =>
					ramrwop <= '0';
					swsrc <= '0';
					aluop <= "0010";
					case if_rf_st(0) is
						when '0' => -- mfih
							dir := "000";
							regwrbop <= "00";
						when '1' => -- mtih
							dir := "110";
							regwrbop <= "00";
						when others =>
							dir := "111";
							regwrbop <= "11";
					end case;
            when others =>
					ramrwop <= '0';
					swsrc <= '0';
					aluop <= "1111";
					dir := "111";
					regwrbop <= "11";
			end case;
			dirop <= dir;
	end process;

	-- ������������չ�Ŀ����ź�
	-- ʹ��IF�εĵõ���IF_INS
    process(IF_Ins)
	-- EX Digits Op
	-- 000 10:0
	-- 001 7:0
	-- 011 4:0
	-- 010 4:2
	-- 110 3:0
	-- others Z... (ILLEGAL)
    begin
        case IF_Ins(15 downto 11) is
            when "01001" => -- addiu
            	ExDigitsOp <= "001";
           		ExSignOp <= '1';
            when "01000" => -- addiu3
            	ExDigitsOp <= "110";
           		ExSignOp <= '1';
            when "01100" => --addsp, bteqz, mtsp
            	if(IF_Ins(10 downto 8)="000" or IF_Ins(10 downto 8)="011") then
            		ExDigitsOp <= "001";
           			ExSignOp <= '1';
           		else
           		end if;
            when "00000" => --addsp3
            	ExDigitsOp <= "001";
           		ExSignOp <= '1';
            when "00010" => -- b
            	ExDigitsOp <= "000";
           		ExSignOp <= '1';
            when "00100" => -- beqz
            	ExDigitsOp <= "001";
           		ExSignOp <= '1';
            when "00101" => -- bnez
            	ExDigitsOp <= "001";
           		ExSignOp <= '1';
            when "01110" => -- cmpi
            	ExDigitsOp <= "001";
           		ExSignOp <= '1';
            when "01101" => -- li
            	ExDigitsOp <= "001";
           		ExSignOp <= '0';
            when "10011" => -- lw
            	ExDigitsOp <= "011";
           		ExSignOp <= '1';
            when "10010" => -- lw_sp
            	ExDigitsOp <= "001";
           		ExSignOp <= '1';
            when "00110" => -- sll, sra
            	ExDigitsOp <= "010";
           		ExSignOp <= '0';
            when "01010" => -- slti
            	ExDigitsOp <= "001";
           		ExSignOp <= '1';
            when "11011" => -- sw
            	ExDigitsOp <= "011";
           		ExSignOp <= '1';
            when "11010" => -- swsp
            	ExDigitsOp <= "001";
           		ExSignOp <= '1';
            when others =>
            	ExDigitsOp <= "111";
           		ExSignOp <= '1';
        end case;
    end process;
    
	 
	-- template
	process
		variable op: STD_LOGIC_VECTOR (4 downto 0);
	begin
		op := if_rf_st (15 downto 11);
		case op is
            when "01001" => -- addiu
            when "01000" => -- addiu3
            when "01100" => 
					case if_rf_st (10 downto 8) is
						when "011" => -- addsp
						when "000" => --btnez
						when "100" => --mtsp
						when others =>
					end case;
            when "00000" => --addsp3
            when "00010" => -- b
            when "00100" => -- beqz
            when "00101" => -- bnez
            when "01110" => -- cmpi
            when "01101" => -- li
            when "10011" => -- lw
            when "10010" => -- lw_sp
            when "00110" => -- sll, sra
					case if_rf_st(1 downto 0) is
						when "00" =>
						when "11" =>
						when others =>
					end case;
            when "01010" => -- slti
				when "01111" => --move
            when "11011" => -- sw
            when "11010" => -- swsp
				when "11100" => 
					case if_rf_st(1 downto 0) is
						when "01" => --addu
						when "11" => --subu
						when others =>
					end case;
				when "11101" =>
					case if_rf_st(4 downto 0) is
						when "01100" => -- add
						when "01010" => --cmp
						when "11101" => --or
						when "00100" => -- sllv
						when "00000" => 
							if if_rf_st(7 downto 5) = "0000" then --jr
							elsif if_rf_st(7 downto 5) = "0100" then --mfpc
							else
							end if;
						when others =>
					end case;
				when "11110" => --mfih and mtih
            when others =>
			end case;
	end process;
end Behavioral;
