----------------------------------------------------------------------------------
-- Company: Concept Computer Corporation
-- Engineer: LXH, LZY, YST
-- 
-- Create Date:    10:29:06 11/19/2016 
-- Design Name: 
-- Module Name:    MemUart - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;

entity MemUart is
    Port ( clk : in STD_LOGIC; --������Ҫ����ʱ��
           rst : in STD_LOGIC; -- ˢ��״̬�� rst='0'����StateΪ00
           
           -- IF
           -- ����PC����ȡָ
           PC_RF_PC : in STD_LOGIC_VECTOR(15 downto 0); --ȡָ��ĵ�ַ
           IF_Ins : out STD_LOGIC_VECTOR(15 downto 0); --ָ�����
           -- MEM
           -- ��ַ��exe_rf_res.
           MEM_SW_DATA : in STD_LOGIC_VECTOR (15 downto 0);
           EXE_RF_Res : in STD_LOGIC_VECTOR(15 downto 0);
           MEM_LW : out STD_LOGIC_VECTOR(15 downto 0);
           
           -- IF & MEM
           -- 0 read; 1 write
           RamRWOp : in std_logic; --�ڴ��д
           
           Addr1 : out STD_LOGIC_VECTOR(15 downto 0);
           Addr2 : out STD_LOGIC_VECTOR(15 downto 0);
           Data1 : inout STD_LOGIC_VECTOR(15 downto 0);  -- low 8 digits for Uart
           Data2 : inout STD_LOGIC_VECTOR(15 downto 0);
           Ram1EN : out STD_LOGIC;
           Ram1OE : out STD_LOGIC;
           Ram1WE : out STD_LOGIC;
           Ram2EN : out STD_LOGIC;
           Ram2OE : out STD_LOGIC;
           Ram2WE : out STD_LOGIC;
           UartRdn : out STD_LOGIC;
           UartWrn : out STD_LOGIC;
			  -------DEBUG--------------
			  state_out : out std_logic_vector (3 downto 0);
           DataReady : in STD_LOGIC;
           Tbre : in STD_LOGIC;
           Tsre : in STD_LOGIC);
end MemUart;

architecture Behavioral of MemUart is
	signal state: STD_LOGIC_VECTOR (1 downto 0) := "00";
	shared variable data : std_logic_vector (15 downto 0) := "0000000000000000";
begin
	state_out <= "00" & state;
	
	process (clk, rst)
		variable write_data : std_logic_vector (15 downto 0) := "0000000000000000";
	begin
		if rst = '0' then
			state <= "00";
		elsif rising_edge (clk) then
			case state is 
				when "00" =>
					if_ins <= "0000100000000000";
					if exe_rf_res(15 downto 2) = "10111111000000" then
						ram1en <= '1';		ram1oe <= '1';		ram1we <= '1';		addr1 <= "ZZZZZZZZZZZZZZZZ";
						ram2en <= '1';		ram2oe <= '1';		ram2we <= '1';		addr2 <= "ZZZZZZZZZZZZZZZZ";
						uartwrn <= '1';	uartrdn <= '1';
						data1 <= "ZZZZZZZZZZZZZZZZ";
						data2 <= "ZZZZZZZZZZZZZZZZ";
					elsif exe_rf_res (15) = '1' then
						ram2en <= '1';		ram2oe <= '1';		ram2we <= '1'; 	addr2 <= "ZZZZZZZZZZZZZZZZ";
						uartwrn <= '1';	uartrdn <= '1';
						data2 <= "ZZZZZZZZZZZZZZZZ";
						if ramrwop = '0' then
							ram1en <= '0';		ram1we <= '1';		ram1oe <= '0';
							data1 <= "ZZZZZZZZZZZZZZZZ";
							addr1 <= exe_rf_res;
						elsif ramrwop = '1' then
							ram1en <= '0';		ram1we <= '1';		ram1oe <= '1';
						else
							ram1en <= '1';		ram1we <= '1';		ram1oe <= '1';
							data1 <= "ZZZZZZZZZZZZZZZZ";
							addr1 <= "ZZZZZZZZZZZZZZZZ";
						end if;
					elsif exe_rf_res(15) = '0' then
						ram1en <= '1';		ram1oe <= '1';		ram1we <= '1';		addr1 <= "ZZZZZZZZZZZZZZZZ";
						uartwrn <= '1';	uartrdn <= '1';
						if ramrwop = '0' then
							ram2en <= '0';		ram2we <= '1';		ram2oe <= '0';
							data2 <= "ZZZZZZZZZZZZZZZZ";
							addr2 <= exe_rf_res;
						elsif ramrwop = '1' then
							ram2en <= '0';		ram2we <= '1';		ram2oe <= '1';
						else
							ram2en <= '1';			ram2we <= '1';		ram2oe <= '1';
							data2 <= "ZZZZZZZZZZZZZZZZ";
							addr2 <= "ZZZZZZZZZZZZZZZZ";
						end if;
					else
						ram1en <= '1';		ram1oe <= '1';		ram1we <= '1';		addr1 <= "ZZZZZZZZZZZZZZZZ";
						ram2en <= '1';		ram2oe <= '1';		ram2we <= '1';	addr2 <= "ZZZZZZZZZZZZZZZZ";
						uartwrn <= '1';	uartrdn <= '1';
					end if;
				when "01" =>
					if exe_rf_res(15 downto 2) = "10111111000000" then
						if ramrwop = '0' then
							uartrdn <= '1';
							uartwrn <= '1';
							data1 <= "ZZZZZZZZZZZZZZZZ";
						elsif ramrwop = '1' then
							data1(7 downto 0) <= mem_sw_data (7 downto 0);
							uartwrn <= '0';
						end if;
					elsif exe_rf_res (15) = '1' then
						if ramrwop = '0' then
							data  := data1;
						elsif ramrwop = '1' then
							data1 <= mem_sw_data;
							ram1we <= '0';
							addr1 <= exe_rf_res;
						end if;
					elsif exe_rf_res(15) = '0' then
						if ramrwop = '0' then
							data := data2;
						elsif ramrwop = '1' then
							data2 <= mem_sw_data;
							ram2we <= '0';
							addr2 <= exe_rf_res;
						end if;
					else
						ram1en <= '1';		ram1oe <= '1';		ram1we <= '1';		addr1 <= "ZZZZZZZZZZZZZZZZ";
						ram2en <= '1';		ram2oe <= '1';		ram2we <= '1';		addr2 <= "ZZZZZZZZZZZZZZZZ";
						uartwrn <= '1';	uartrdn <= '1';
					end if;
				when "10" =>
					ram1en <= '1';		ram1oe <= '1';		ram1we <= '1';
					if exe_rf_res(15 downto 2) = "10111111000000" then
						if ramrwop = '0' then
							uartwrn <= '1';
							uartrdn <= '0';
						else
							uartwrn <= '1';
						end if;
					end if;
					ram2en <= '0';	ram2oe <= '0';	ram2we <= '1';
					data2 <= "ZZZZZZZZZZZZZZZZ";
					addr2 <= pc_rf_pc;
				when "11" =>
					if exe_rf_res(15 downto 2) = "10111111000000" then
						if ramrwop = '0' then
							if exe_rf_res(0) = '0' then
								data := "00000000" & data1(7 downto 0);
							else
								data := "00000000000000" & dataready & (tbre and tsre);
							end if;
						end if;
					end if;
					if_ins <= data2;
				when others =>
					if_ins <= "0000100000000000";
					data := "1111111111111111";
					addr1 <= "ZZZZZZZZZZZZZZZZ";
					addr2 <= "ZZZZZZZZZZZZZZZZ";
					ram1en <= '1';
					ram1we <= '1';
					ram1oe <= '1';
					ram2en <= '1';
					ram2oe <= '1';
					ram2we <= '1';
					uartwrn <= '1';
					uartrdn <= '1';
			end case;
			mem_lw <= data;
			state <= state + 1;
		end if;
	end process;
end Behavioral;
